// ------------
// SPI RTL-code header

`include "fifo.v"
`include "baud_rate_gen.v"
`include "spi_transceiver.v"
`include "spi_control.v"
`include "spi_top.v"

// ------------
